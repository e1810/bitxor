module AND(
	input wire in0,
	input wire in1,
	output wire out0
	);

	assign out0 = in0 & in1;
endmodule
